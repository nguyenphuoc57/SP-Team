module int2float (in, out);

input [7:0] in;
output reg [31:0] out;

always @(in) begin
	case(in) 
	8'h00: out = 32'h0;
        8'h01: out = 32'h3b808081;
        8'h02: out = 32'h3c008081;
        8'h03: out = 32'h3c40c0c1;
        8'h04: out = 32'h3c808081;
        8'h05: out = 32'h3ca0a0a1;
        8'h06: out = 32'h3cc0c0c1;
        8'h07: out = 32'h3ce0e0e1;
        8'h08: out = 32'h3d008081;
        8'h09: out = 32'h3d109091;
        8'h0a: out = 32'h3d20a0a1;
        8'h0b: out = 32'h3d30b0b1;
        8'h0c: out = 32'h3d40c0c1;
        8'h0d: out = 32'h3d50d0d1;
        8'h0e: out = 32'h3d60e0e1;
        8'h0f: out = 32'h3d70f0f1;
        8'h10: out = 32'h3d808081;
        8'h11: out = 32'h3d888889;
        8'h12: out = 32'h3d909091;
        8'h13: out = 32'h3d989899;
        8'h14: out = 32'h3da0a0a1;
        8'h15: out = 32'h3da8a8a9;
        8'h16: out = 32'h3db0b0b1;
        8'h17: out = 32'h3db8b8b9;
        8'h18: out = 32'h3dc0c0c1;
        8'h19: out = 32'h3dc8c8c9;
        8'h1a: out = 32'h3dd0d0d1;
        8'h1b: out = 32'h3dd8d8d9;
        8'h1c: out = 32'h3de0e0e1;
        8'h1d: out = 32'h3de8e8e9;
        8'h1e: out = 32'h3df0f0f1;
        8'h1f: out = 32'h3df8f8f9;
        8'h20: out = 32'h3e008081;
        8'h21: out = 32'h3e048485;
        8'h22: out = 32'h3e088889;
        8'h23: out = 32'h3e0c8c8d;
        8'h24: out = 32'h3e109091;
        8'h25: out = 32'h3e149495;
        8'h26: out = 32'h3e189899;
        8'h27: out = 32'h3e1c9c9d;
        8'h28: out = 32'h3e20a0a1;
        8'h29: out = 32'h3e24a4a5;
        8'h2a: out = 32'h3e28a8a9;
        8'h2b: out = 32'h3e2cacad;
        8'h2c: out = 32'h3e30b0b1;
        8'h2d: out = 32'h3e34b4b5;
        8'h2e: out = 32'h3e38b8b9;
        8'h2f: out = 32'h3e3cbcbd;
        8'h30: out = 32'h3e40c0c1;
        8'h31: out = 32'h3e44c4c5;
        8'h32: out = 32'h3e48c8c9;
        8'h33: out = 32'h3e4ccccd;
        8'h34: out = 32'h3e50d0d1;
        8'h35: out = 32'h3e54d4d5;
        8'h36: out = 32'h3e58d8d9;
        8'h37: out = 32'h3e5cdcdd;
        8'h38: out = 32'h3e60e0e1;
        8'h39: out = 32'h3e64e4e5;
        8'h3a: out = 32'h3e68e8e9;
        8'h3b: out = 32'h3e6ceced;
        8'h3c: out = 32'h3e70f0f1;
        8'h3d: out = 32'h3e74f4f5;
        8'h3e: out = 32'h3e78f8f9;
        8'h3f: out = 32'h3e7cfcfd;
        8'h40: out = 32'h3e808081;
        8'h41: out = 32'h3e828283;
        8'h42: out = 32'h3e848485;
        8'h43: out = 32'h3e868687;
        8'h44: out = 32'h3e888889;
        8'h45: out = 32'h3e8a8a8b;
        8'h46: out = 32'h3e8c8c8d;
        8'h47: out = 32'h3e8e8e8f;
        8'h48: out = 32'h3e909091;
        8'h49: out = 32'h3e929293;
        8'h4a: out = 32'h3e949495;
        8'h4b: out = 32'h3e969697;
        8'h4c: out = 32'h3e989899;
        8'h4d: out = 32'h3e9a9a9b;
        8'h4e: out = 32'h3e9c9c9d;
        8'h4f: out = 32'h3e9e9e9f;
        8'h50: out = 32'h3ea0a0a1;
        8'h51: out = 32'h3ea2a2a3;
        8'h52: out = 32'h3ea4a4a5;
        8'h53: out = 32'h3ea6a6a7;
        8'h54: out = 32'h3ea8a8a9;
        8'h55: out = 32'h3eaaaaab;
        8'h56: out = 32'h3eacacad;
        8'h57: out = 32'h3eaeaeaf;
        8'h58: out = 32'h3eb0b0b1;
        8'h59: out = 32'h3eb2b2b3;
        8'h5a: out = 32'h3eb4b4b5;
        8'h5b: out = 32'h3eb6b6b7;
        8'h5c: out = 32'h3eb8b8b9;
        8'h5d: out = 32'h3ebababb;
        8'h5e: out = 32'h3ebcbcbd;
        8'h5f: out = 32'h3ebebebf;
        8'h60: out = 32'h3ec0c0c1;
        8'h61: out = 32'h3ec2c2c3;
        8'h62: out = 32'h3ec4c4c5;
        8'h63: out = 32'h3ec6c6c7;
        8'h64: out = 32'h3ec8c8c9;
        8'h65: out = 32'h3ecacacb;
        8'h66: out = 32'h3ecccccd;
        8'h67: out = 32'h3ecececf;
        8'h68: out = 32'h3ed0d0d1;
        8'h69: out = 32'h3ed2d2d3;
        8'h6a: out = 32'h3ed4d4d5;
        8'h6b: out = 32'h3ed6d6d7;
        8'h6c: out = 32'h3ed8d8d9;
        8'h6d: out = 32'h3edadadb;
        8'h6e: out = 32'h3edcdcdd;
        8'h6f: out = 32'h3edededf;
        8'h70: out = 32'h3ee0e0e1;
        8'h71: out = 32'h3ee2e2e3;
        8'h72: out = 32'h3ee4e4e5;
        8'h73: out = 32'h3ee6e6e7;
        8'h74: out = 32'h3ee8e8e9;
        8'h75: out = 32'h3eeaeaeb;
        8'h76: out = 32'h3eececed;
        8'h77: out = 32'h3eeeeeef;
        8'h78: out = 32'h3ef0f0f1;
        8'h79: out = 32'h3ef2f2f3;
        8'h7a: out = 32'h3ef4f4f5;
        8'h7b: out = 32'h3ef6f6f7;
        8'h7c: out = 32'h3ef8f8f9;
        8'h7d: out = 32'h3efafafb;
        8'h7e: out = 32'h3efcfcfd;
        8'h7f: out = 32'h3efefeff;
        8'h80: out = 32'h3f008081;
        8'h81: out = 32'h3f018182;
        8'h82: out = 32'h3f028283;
        8'h83: out = 32'h3f038384;
        8'h84: out = 32'h3f048485;
        8'h85: out = 32'h3f058586;
        8'h86: out = 32'h3f068687;
        8'h87: out = 32'h3f078788;
        8'h88: out = 32'h3f088889;
        8'h89: out = 32'h3f09898a;
        8'h8a: out = 32'h3f0a8a8b;
        8'h8b: out = 32'h3f0b8b8c;
        8'h8c: out = 32'h3f0c8c8d;
        8'h8d: out = 32'h3f0d8d8e;
        8'h8e: out = 32'h3f0e8e8f;
        8'h8f: out = 32'h3f0f8f90;
        8'h90: out = 32'h3f109091;
        8'h91: out = 32'h3f119192;
        8'h92: out = 32'h3f129293;
        8'h93: out = 32'h3f139394;
        8'h94: out = 32'h3f149495;
        8'h95: out = 32'h3f159596;
        8'h96: out = 32'h3f169697;
        8'h97: out = 32'h3f179798;
        8'h98: out = 32'h3f189899;
        8'h99: out = 32'h3f19999a;
        8'h9a: out = 32'h3f1a9a9b;
        8'h9b: out = 32'h3f1b9b9c;
        8'h9c: out = 32'h3f1c9c9d;
        8'h9d: out = 32'h3f1d9d9e;
        8'h9e: out = 32'h3f1e9e9f;
        8'h9f: out = 32'h3f1f9fa0;
        8'ha0: out = 32'h3f20a0a1;
        8'ha1: out = 32'h3f21a1a2;
        8'ha2: out = 32'h3f22a2a3;
        8'ha3: out = 32'h3f23a3a4;
        8'ha4: out = 32'h3f24a4a5;
        8'ha5: out = 32'h3f25a5a6;
        8'ha6: out = 32'h3f26a6a7;
        8'ha7: out = 32'h3f27a7a8;
        8'ha8: out = 32'h3f28a8a9;
        8'ha9: out = 32'h3f29a9aa;
        8'haa: out = 32'h3f2aaaab;
        8'hab: out = 32'h3f2babac;
        8'hac: out = 32'h3f2cacad;
        8'had: out = 32'h3f2dadae;
        8'hae: out = 32'h3f2eaeaf;
        8'haf: out = 32'h3f2fafb0;
        8'hb0: out = 32'h3f30b0b1;
        8'hb1: out = 32'h3f31b1b2;
        8'hb2: out = 32'h3f32b2b3;
        8'hb3: out = 32'h3f33b3b4;
        8'hb4: out = 32'h3f34b4b5;
        8'hb5: out = 32'h3f35b5b6;
        8'hb6: out = 32'h3f36b6b7;
        8'hb7: out = 32'h3f37b7b8;
        8'hb8: out = 32'h3f38b8b9;
        8'hb9: out = 32'h3f39b9ba;
        8'hba: out = 32'h3f3ababb;
        8'hbb: out = 32'h3f3bbbbc;
        8'hbc: out = 32'h3f3cbcbd;
        8'hbd: out = 32'h3f3dbdbe;
        8'hbe: out = 32'h3f3ebebf;
        8'hbf: out = 32'h3f3fbfc0;
        8'hc0: out = 32'h3f40c0c1;
        8'hc1: out = 32'h3f41c1c2;
        8'hc2: out = 32'h3f42c2c3;
        8'hc3: out = 32'h3f43c3c4;
        8'hc4: out = 32'h3f44c4c5;
        8'hc5: out = 32'h3f45c5c6;
        8'hc6: out = 32'h3f46c6c7;
        8'hc7: out = 32'h3f47c7c8;
        8'hc8: out = 32'h3f48c8c9;
        8'hc9: out = 32'h3f49c9ca;
        8'hca: out = 32'h3f4acacb;
        8'hcb: out = 32'h3f4bcbcc;
        8'hcc: out = 32'h3f4ccccd;
        8'hcd: out = 32'h3f4dcdce;
        8'hce: out = 32'h3f4ececf;
        8'hcf: out = 32'h3f4fcfd0;
        8'hd0: out = 32'h3f50d0d1;
        8'hd1: out = 32'h3f51d1d2;
        8'hd2: out = 32'h3f52d2d3;
        8'hd3: out = 32'h3f53d3d4;
        8'hd4: out = 32'h3f54d4d5;
        8'hd5: out = 32'h3f55d5d6;
        8'hd6: out = 32'h3f56d6d7;
        8'hd7: out = 32'h3f57d7d8;
        8'hd8: out = 32'h3f58d8d9;
        8'hd9: out = 32'h3f59d9da;
        8'hda: out = 32'h3f5adadb;
        8'hdb: out = 32'h3f5bdbdc;
        8'hdc: out = 32'h3f5cdcdd;
        8'hdd: out = 32'h3f5dddde;
        8'hde: out = 32'h3f5ededf;
        8'hdf: out = 32'h3f5fdfe0;
        8'he0: out = 32'h3f60e0e1;
        8'he1: out = 32'h3f61e1e2;
        8'he2: out = 32'h3f62e2e3;
        8'he3: out = 32'h3f63e3e4;
        8'he4: out = 32'h3f64e4e5;
        8'he5: out = 32'h3f65e5e6;
        8'he6: out = 32'h3f66e6e7;
        8'he7: out = 32'h3f67e7e8;
        8'he8: out = 32'h3f68e8e9;
        8'he9: out = 32'h3f69e9ea;
        8'hea: out = 32'h3f6aeaeb;
        8'heb: out = 32'h3f6bebec;
        8'hec: out = 32'h3f6ceced;
        8'hed: out = 32'h3f6dedee;
        8'hee: out = 32'h3f6eeeef;
        8'hef: out = 32'h3f6feff0;
        8'hf0: out = 32'h3f70f0f1;
        8'hf1: out = 32'h3f71f1f2;
        8'hf2: out = 32'h3f72f2f3;
        8'hf3: out = 32'h3f73f3f4;
        8'hf4: out = 32'h3f74f4f5;
        8'hf5: out = 32'h3f75f5f6;
        8'hf6: out = 32'h3f76f6f7;
        8'hf7: out = 32'h3f77f7f8;
        8'hf8: out = 32'h3f78f8f9;
        8'hf9: out = 32'h3f79f9fa;
        8'hfa: out = 32'h3f7afafb;
	8'hfb: out = 32'h3f7bfbfc;
        8'hfc: out = 32'h3f7cfcfd;
        8'hfd: out = 32'h3f7dfdfe;
        8'hfe: out = 32'h3f7efeff;
        8'hff: out = 32'h3F800000;
	default: out=32'h0;
endcase
end
endmodule
module layer1 (clk,reset,enable_conv,enable_max,data_in_1, 
data_in_2, 
data_in_3, 
data_in_4, 
data_in_5, 
data_in_6, 
data_in_7, 
data_in_8, 
data_in_9, 
data_in_10, 
data_in_11, 
data_in_12, 
data_in_13, 
data_in_14, 
data_in_15, 
data_in_16, 
data_in_17, 
data_in_18, 
data_in_19, 
data_in_20, 
data_in_21, 
data_in_22, 
data_in_23, 
data_in_24, 
data_in_25, 
data_in_26, 
data_in_27, 
data_in_28, 
data_in_29, 
data_in_30, 
data_in_31, 
data_in_32, 
data_in_33, 
data_in_34, 
data_in_35, 
data_in_36, 
data_in_37, 
data_in_38, 
data_in_39, 
data_in_40, 
data_in_41, 
data_in_42, 
data_in_43, 
data_in_44, 
data_in_45, 
data_in_46, 
data_in_47, 
data_in_48, 
data_in_49, 
data_in_50, 
data_in_51, 
data_in_52, 
data_in_53, 
data_in_54, 
data_in_55, 
data_in_56, 
data_in_57, 
data_in_58, 
data_in_59, 
data_in_60, 
data_in_61, 
data_in_62, 
data_in_63, 
data_in_64, 
	kernel_in_1,
	kernel_in_2,
	kernel_in_3,
	kernel_in_4,
	kernel_in_5,
	kernel_in_6,
	kernel_in_7,
	kernel_in_8,
	kernel_in_9,
	kernel_in_10,
	kernel_in_11,
	kernel_in_12,
	kernel_in_13,
	kernel_in_14,
	kernel_in_15,
	kernel_in_16,
	kernel_in_17,
	kernel_in_18,
	kernel_in_19,
	kernel_in_20,
	kernel_in_21,
	kernel_in_22,
	kernel_in_23,
	kernel_in_24,
	kernel_in_25,
	kernel_in_26,
	kernel_in_27,
	kernel_in_28,
	kernel_in_29,
	kernel_in_30,
	kernel_in_31,
	kernel_in_32,
	kernel_in_33,
	kernel_in_34,
	kernel_in_35,
	kernel_in_36,
	kernel_in_37,
	kernel_in_38,
	kernel_in_39,
	kernel_in_40,
	kernel_in_41,
	kernel_in_42,
	kernel_in_43,
	kernel_in_44,
	kernel_in_45,
	kernel_in_46,
	kernel_in_47,
	kernel_in_48,
	kernel_in_49,
	kernel_in_50,
	kernel_in_51,
	kernel_in_52,
	kernel_in_53,
	kernel_in_54,
	kernel_in_55,
	kernel_in_56,
	kernel_in_57,
	kernel_in_58,
	kernel_in_59,
	kernel_in_60,
	kernel_in_61,
	kernel_in_62,
	kernel_in_63,
	kernel_in_64,
	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	data_out_9,
	data_out_10,
	data_out_11,
	data_out_12,
	data_out_13,
	data_out_14,
	data_out_15,
	data_out_16,
	data_out_17,
	data_out_18,
	data_out_19,
	data_out_20,
	data_out_21,
	data_out_22,
	data_out_23,
	data_out_24,
	data_out_25,
	data_out_26,
	data_out_27,
	data_out_28,
	data_out_29,
	data_out_30,
	data_out_31,
	data_out_32,
	data_out_33,
	data_out_34,
	data_out_35,
	data_out_36,
	data_out_37,
	data_out_38,
	data_out_39,
	data_out_40,
	data_out_41,
	data_out_42,
	data_out_43,
	data_out_44,
	data_out_45,
	data_out_46,
	data_out_47,
	data_out_48,
	data_out_49,
	data_out_50,
	data_out_51,
	data_out_52,
	data_out_53,
	data_out_54,
	data_out_55,
	data_out_56,
	data_out_57,
	data_out_58,
	data_out_59,
	data_out_60,
	data_out_61,
	data_out_62,
	data_out_63,
	data_out_64,
valid_in, valid_out
);
input clk,reset,enable_conv, enable_max;
input [31:0] 		data_in_1, 
		data_in_2, 
		data_in_3, 
		data_in_4, 
		data_in_5, 
		data_in_6, 
		data_in_7, 
		data_in_8, 
		data_in_9, 
		data_in_10, 
		data_in_11, 
		data_in_12, 
		data_in_13, 
		data_in_14, 
		data_in_15, 
		data_in_16, 
		data_in_17, 
		data_in_18, 
		data_in_19, 
		data_in_20, 
		data_in_21, 
		data_in_22, 
		data_in_23, 
		data_in_24, 
		data_in_25, 
		data_in_26, 
		data_in_27, 
		data_in_28, 
		data_in_29, 
		data_in_30, 
		data_in_31, 
		data_in_32, 
		data_in_33, 
		data_in_34, 
		data_in_35, 
		data_in_36, 
		data_in_37, 
		data_in_38, 
		data_in_39, 
		data_in_40, 
		data_in_41, 
		data_in_42, 
		data_in_43, 
		data_in_44, 
		data_in_45, 
		data_in_46, 
		data_in_47, 
		data_in_48, 
		data_in_49, 
		data_in_50, 
		data_in_51, 
		data_in_52, 
		data_in_53, 
		data_in_54, 
		data_in_55, 
		data_in_56, 
		data_in_57, 
		data_in_58, 
		data_in_59, 
		data_in_60, 
		data_in_61, 
		data_in_62, 
		data_in_63, 
		data_in_64, 
		kernel_in_1,
		kernel_in_2,
		kernel_in_3,
		kernel_in_4,
		kernel_in_5,
		kernel_in_6,
		kernel_in_7,
		kernel_in_8,
		kernel_in_9,
		kernel_in_10,
		kernel_in_11,
		kernel_in_12,
		kernel_in_13,
		kernel_in_14,
		kernel_in_15,
		kernel_in_16,
		kernel_in_17,
		kernel_in_18,
		kernel_in_19,
		kernel_in_20,
		kernel_in_21,
		kernel_in_22,
		kernel_in_23,
		kernel_in_24,
		kernel_in_25,
		kernel_in_26,
		kernel_in_27,
		kernel_in_28,
		kernel_in_29,
		kernel_in_30,
		kernel_in_31,
		kernel_in_32,
		kernel_in_33,
		kernel_in_34,
		kernel_in_35,
		kernel_in_36,
		kernel_in_37,
		kernel_in_38,
		kernel_in_39,
		kernel_in_40,
		kernel_in_41,
		kernel_in_42,
		kernel_in_43,
		kernel_in_44,
		kernel_in_45,
		kernel_in_46,
		kernel_in_47,
		kernel_in_48,
		kernel_in_49,
		kernel_in_50,
		kernel_in_51,
		kernel_in_52,
		kernel_in_53,
		kernel_in_54,
		kernel_in_55,
		kernel_in_56,
		kernel_in_57,
		kernel_in_58,
		kernel_in_59,
		kernel_in_60,
		kernel_in_61,
		kernel_in_62,
		kernel_in_63,
		kernel_in_64,
;
output valid_in, valid_out; 
output [31:0] 	data_out_1,
	data_out_2,
	data_out_3,
	data_out_4,
	data_out_5,
	data_out_6,
	data_out_7,
	data_out_8,
	data_out_9,
	data_out_10,
	data_out_11,
	data_out_12,
	data_out_13,
	data_out_14,
	data_out_15,
	data_out_16,
	data_out_17,
	data_out_18,
	data_out_19,
	data_out_20,
	data_out_21,
	data_out_22,
	data_out_23,
	data_out_24,
	data_out_25,
	data_out_26,
	data_out_27,
	data_out_28,
	data_out_29,
	data_out_30,
	data_out_31,
	data_out_32,
	data_out_33,
	data_out_34,
	data_out_35,
	data_out_36,
	data_out_37,
	data_out_38,
	data_out_39,
	data_out_40,
	data_out_41,
	data_out_42,
	data_out_43,
	data_out_44,
	data_out_45,
	data_out_46,
	data_out_47,
	data_out_48,
	data_out_49,
	data_out_50,
	data_out_51,
	data_out_52,
	data_out_53,
	data_out_54,
	data_out_55,
	data_out_56,
	data_out_57,
	data_out_58,
	data_out_59,
	data_out_60,
	data_out_61,
	data_out_62,
	data_out_63,
	data_out_64,
block1 1( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_1),
		   .kernel_in(kernel_in_1),
		   .data_out(data_out_1),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 2( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_2),
		   .kernel_in(kernel_in_2),
		   .data_out(data_out_2),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 3( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_3),
		   .kernel_in(kernel_in_3),
		   .data_out(data_out_3),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 4( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_4),
		   .kernel_in(kernel_in_4),
		   .data_out(data_out_4),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 5( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_5),
		   .kernel_in(kernel_in_5),
		   .data_out(data_out_5),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 6( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_6),
		   .kernel_in(kernel_in_6),
		   .data_out(data_out_6),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 7( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_7),
		   .kernel_in(kernel_in_7),
		   .data_out(data_out_7),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 8( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_8),
		   .kernel_in(kernel_in_8),
		   .data_out(data_out_8),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 9( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_9),
		   .kernel_in(kernel_in_9),
		   .data_out(data_out_9),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 10( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_10),
		   .kernel_in(kernel_in_10),
		   .data_out(data_out_10),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 11( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_11),
		   .kernel_in(kernel_in_11),
		   .data_out(data_out_11),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 12( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_12),
		   .kernel_in(kernel_in_12),
		   .data_out(data_out_12),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 13( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_13),
		   .kernel_in(kernel_in_13),
		   .data_out(data_out_13),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 14( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_14),
		   .kernel_in(kernel_in_14),
		   .data_out(data_out_14),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 15( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_15),
		   .kernel_in(kernel_in_15),
		   .data_out(data_out_15),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 16( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_16),
		   .kernel_in(kernel_in_16),
		   .data_out(data_out_16),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 17( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_17),
		   .kernel_in(kernel_in_17),
		   .data_out(data_out_17),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 18( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_18),
		   .kernel_in(kernel_in_18),
		   .data_out(data_out_18),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 19( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_19),
		   .kernel_in(kernel_in_19),
		   .data_out(data_out_19),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 20( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_20),
		   .kernel_in(kernel_in_20),
		   .data_out(data_out_20),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 21( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_21),
		   .kernel_in(kernel_in_21),
		   .data_out(data_out_21),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 22( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_22),
		   .kernel_in(kernel_in_22),
		   .data_out(data_out_22),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 23( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_23),
		   .kernel_in(kernel_in_23),
		   .data_out(data_out_23),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 24( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_24),
		   .kernel_in(kernel_in_24),
		   .data_out(data_out_24),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 25( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_25),
		   .kernel_in(kernel_in_25),
		   .data_out(data_out_25),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 26( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_26),
		   .kernel_in(kernel_in_26),
		   .data_out(data_out_26),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 27( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_27),
		   .kernel_in(kernel_in_27),
		   .data_out(data_out_27),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 28( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_28),
		   .kernel_in(kernel_in_28),
		   .data_out(data_out_28),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 29( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_29),
		   .kernel_in(kernel_in_29),
		   .data_out(data_out_29),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 30( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_30),
		   .kernel_in(kernel_in_30),
		   .data_out(data_out_30),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 31( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_31),
		   .kernel_in(kernel_in_31),
		   .data_out(data_out_31),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 32( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_32),
		   .kernel_in(kernel_in_32),
		   .data_out(data_out_32),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 33( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_33),
		   .kernel_in(kernel_in_33),
		   .data_out(data_out_33),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 34( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_34),
		   .kernel_in(kernel_in_34),
		   .data_out(data_out_34),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 35( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_35),
		   .kernel_in(kernel_in_35),
		   .data_out(data_out_35),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 36( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_36),
		   .kernel_in(kernel_in_36),
		   .data_out(data_out_36),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 37( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_37),
		   .kernel_in(kernel_in_37),
		   .data_out(data_out_37),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 38( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_38),
		   .kernel_in(kernel_in_38),
		   .data_out(data_out_38),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 39( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_39),
		   .kernel_in(kernel_in_39),
		   .data_out(data_out_39),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 40( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_40),
		   .kernel_in(kernel_in_40),
		   .data_out(data_out_40),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 41( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_41),
		   .kernel_in(kernel_in_41),
		   .data_out(data_out_41),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 42( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_42),
		   .kernel_in(kernel_in_42),
		   .data_out(data_out_42),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 43( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_43),
		   .kernel_in(kernel_in_43),
		   .data_out(data_out_43),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 44( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_44),
		   .kernel_in(kernel_in_44),
		   .data_out(data_out_44),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 45( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_45),
		   .kernel_in(kernel_in_45),
		   .data_out(data_out_45),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 46( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_46),
		   .kernel_in(kernel_in_46),
		   .data_out(data_out_46),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 47( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_47),
		   .kernel_in(kernel_in_47),
		   .data_out(data_out_47),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 48( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_48),
		   .kernel_in(kernel_in_48),
		   .data_out(data_out_48),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 49( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_49),
		   .kernel_in(kernel_in_49),
		   .data_out(data_out_49),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 50( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_50),
		   .kernel_in(kernel_in_50),
		   .data_out(data_out_50),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 51( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_51),
		   .kernel_in(kernel_in_51),
		   .data_out(data_out_51),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 52( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_52),
		   .kernel_in(kernel_in_52),
		   .data_out(data_out_52),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 53( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_53),
		   .kernel_in(kernel_in_53),
		   .data_out(data_out_53),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 54( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_54),
		   .kernel_in(kernel_in_54),
		   .data_out(data_out_54),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 55( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_55),
		   .kernel_in(kernel_in_55),
		   .data_out(data_out_55),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 56( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_56),
		   .kernel_in(kernel_in_56),
		   .data_out(data_out_56),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 57( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_57),
		   .kernel_in(kernel_in_57),
		   .data_out(data_out_57),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 58( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_58),
		   .kernel_in(kernel_in_58),
		   .data_out(data_out_58),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 59( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_59),
		   .kernel_in(kernel_in_59),
		   .data_out(data_out_59),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 60( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_60),
		   .kernel_in(kernel_in_60),
		   .data_out(data_out_60),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 61( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_61),
		   .kernel_in(kernel_in_61),
		   .data_out(data_out_61),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 62( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_62),
		   .kernel_in(kernel_in_62),
		   .data_out(data_out_62),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 63( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_63),
		   .kernel_in(kernel_in_63),
		   .data_out(data_out_63),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
block1 64( .clk(clk),
		   .reset(reset),
		   .enable_conv(enable_conv),
		   .enable_max(enable_max),
		   .data_in(data_in_64),
		   .kernel_in(kernel_in_64),
		   .data_out(data_out_64),
		   .valid_in(valid_in),
		   .valid_out(valid_out)
	);
endmodule

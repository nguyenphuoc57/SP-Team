module fp_add (A,B,C,enable, clk);
input clk;
input [31:0] A,B;
input enable;
output reg [31:0] C;

reg [23:0] ManA, ManB;
reg [24:0] C1;
reg[7:0] expTemp;
reg [24:0] ManC;
reg [7:0] ea, eb;

always @(negedge clk) begin
if (!enable) begin
	C=32'b0;
	ManA = 0;
	ManB=0;
	ea=0;
	eb=0;
end 
else if (A==32'b0 && B==32'b0) begin
	C=32'b0;
end
else begin 
			ManA = {1'd1,A[22:0]};
			ManB= {1'd1,B[22:0]};
			ea= A[30:23];
			eb=B[30:23];	
if (ea< eb) begin     		// A'exp < B'exp
		expTemp = eb - ea;
		ea = eb;
		ManA = ManA >> expTemp;
end 
else begin 											//A'exp >=  B'exp
		expTemp= ea - eb;
		eb = ea;
		ManB = ManB >> expTemp;
end 

if (A[31]==B[31]) begin
	ManC=ManB + ManA;
   C[31] = A[31];
end
else 	if(ManA > ManB) begin 			   // A > B
				ManC= ManA-ManB;
				C[31]=A[31];
			end
else if (ManA < ManB) begin			// A < B
				ManC=ManB - ManA;
				C[31]=B[31];
				end
else begin			// A = B	
					ManC = ManA-ManB;
					C[31] = 1'd0;
				end

if (ManC[24]==1) begin		
				C[22:0]=ManC[23:1];
				C[30:23]=ea+8'd1;
		end
		else if(ManC[23]==1) begin 					
				C[22:0]=ManC[22:0];
				C[30:23]=ea;
		end
		else if (ManC[22]==1) begin
					C[22:0]={ManC[21:0],1'd0};
					C[30:23]=ea-8'd1;
				end
		else if (ManC[21]==1) begin
					C[22:0]={ManC[20:0],2'd0};
					C[30:23]=ea-8'd2;	
				end
		else if (ManC[20]==1) begin
					C[22:0]={ManC[19:0],3'd0};
					C[30:23]=ea-8'd3;	
				end
		else if (ManC[19]==1) begin
					C[22:0]={ManC[18:0],4'd0};
					C[30:23]=ea-8'd4;
				end
		else if (ManC[18]==1) begin
					C[22:0]={ManC[17:0],5'd0};
					C[30:23]=ea-8'd5;
				end
		else if (ManC[17]==1) begin
					C[22:0]={ManC[16:0],6'd0};
					C[30:23]=ea-8'd6;
				end		
		else if (ManC[16]==1) begin
					C[22:0]={ManC[15:0],7'd0};
					C[30:23]=ea-8'd7;
				end		
		else if (ManC[15]==1) begin
					C[22:0]={ManC[14:0],8'd0};
					C[30:23]=ea-8'd8;
				end
		else if (ManC[14]==1) begin
					C[22:0]={ManC[13:0],9'd0};
					C[30:23]=ea-8'd9;
				end
		else if (ManC[13]==1) begin
					C[22:0]={ManC[12:0],10'd0};
					C[30:23]=ea-8'd10;
				end
		else if (ManC[12]==1) begin
					C[22:0]={ManC[11:0],11'd0};
					C[30:23]=ea-8'd11;
				end
		else if (ManC[11]==1) begin
					C[22:0]={ManC[10:0],12'd0};
					C[30:23]=ea-8'd12;
				end
		else if (ManC[10]==1) begin
					C[22:0]={ManC[9:0],13'd0};
					C[30:23]=ea-8'd13;
				end
		else if (ManC[9]==1) begin
					C[22:0]={ManC[8:0],14'd0};
					C[30:23]=ea-8'd14;
				end
		else if (ManC[8]==1) begin
					C[22:0]={ManC[7:0],15'd0};
					C[30:23]=ea-8'd15;
				end
		else if (ManC[7]==1) begin
					C[22:0]={ManC[6:0],16'd0};
					C[30:23]=ea-8'd16;
				end
		else if (ManC[6]==1) begin
					C[22:0]={ManC[5:0],17'd0};
					C[30:23]=ea-8'd17;
				end
		else if (ManC[5]==1) begin
					C[22:0]={ManC[4:0],18'd0};
					C[30:23]=ea-8'd18;
				end
		else if (ManC[4]==1) begin
					C[22:0]={ManC[3:0],19'd0};
					C[30:23]=ea-8'd19;
				end
		else if (ManC[3]==1) begin
					C[22:0]={ManC[2:0],20'd0};
					C[30:23]=ea-8'd20;
				end
		else if (ManC[2]==1) begin
					C[22:0]={ManC[1:0],21'd0};
					C[30:23]=ea-8'd21;
				end
		else if (ManC[1]==1) begin
					C[22:0]={ManC[0],22'd0};
					C[30:23]=ea-8'd22;
				end
		else if (ManC[0]==1) begin
					C[22:0]={23'd0};
					C[30:23]=ea-8'd23;
				end
		else C[30:0]=31'b0;			
end
end
endmodule 

